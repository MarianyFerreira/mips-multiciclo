library ieee;
use ieee.std_logic_1164.all;

entity toplevel is
	port( 	input	: in std_logic_vector (31 downto 0);

				output : out std_logic_vector (31 downto 0)
	);
end ;

architecture arch of toplevel is
	
	-- signal
	
	begin	
	end arch;
