library ieee;
use ieee.std_logic_1164.all;

entity name is
	port( sel : in std_logic_vector (1 downto 0);
			input : in std_logic_vector(31 downto 0);
        	
        	output : out std_logic_vector(31 downto 0)
    );
end;

architecture behavior of name is
	begin
	end behavior;