library ieee;
use ieee.std_logic_1164.all;

entity  nome is
port (
	 );
end  nome ;

architecture arch of  nome  is

	signal
	
	begin
	
	end arch;
